`timescale 1ns / 1ps
module RAM_B (
input wire clka,
input wire wea, 
input wire [5:0] addra,
input wire [31:0] dina, 
output wire [31:0] douta 
);



endmodule
